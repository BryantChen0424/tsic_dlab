module minmax (
    
);
    always @(*) begin
        /* assignment */
    end
endmodule
