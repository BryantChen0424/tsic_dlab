module between (
    
);
    always @(*) begin
        /* assignment */
    end
endmodule
