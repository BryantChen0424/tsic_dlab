module math (
    
);
    always @(*) begin
        
    end
endmodule
