module ops (
    
);

    always @(*) begin

    end
endmodule
