module mul (
    
);
    always @(*) begin
        /* */
    end
endmodule
