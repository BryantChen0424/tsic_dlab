module between (
    input  [7:0] a,
    output reg bt // = if 25 < a < 125 ? 1 for yes, 0 for no.
);
    always @(*) begin
        bt = //
    end
endmodule
